module muxFive(m_out,A,B,select);  
output [4:0] m_out;  input [4:0] A,B;  input select; 
 
 assign m_out = (select)? B:A; 

endmodule 
